library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity Servos is port(
	SX : out std_logic_vector (1 downto 0);
	SY : out std_logic_vector (1 downto 0);
	s1 : out std_logic;
	s2 : out std_logic;
	clock : in std_logic;
	VRX : in std_logic_vector(9 downto 0);
	VRY : in std_logic_vector(9 downto 0));
end Servos;

architecture Behavioral of Servos is 
	signal clk,clktope,relogio,uhr,T,mov0,mov1,mov2: std_logic := '1';
	signal cont,cont1,cont0 : integer := 1;
	signal s�0,s�1,s�2,s�3,s�4,s�5,s�6,s�7,s�8,s�9,s�10 : std_logic := '1';
	signal s�11,s�12,s�13,s�14,s�15,s�16,s�17,s�18,s�19 : std_logic := '1';
	signal se�al : std_logic_vector (5 downto 0) := "000001";
	signal doscientos: std_logic_vector (7 downto 0) := "00000001";
	signal se�alt : std_logic_vector (4 downto 0) := "00001";
begin
clk <= clock;

--------------------Main Process-----------------------
	process (VRY, VRX, mov0, mov1, mov2, relogio) begin
	---Parte Servomotor con 360� de libertad
		if VRY < "0100101100" then
			SY <= "01";
			s1 <= mov1;
		elsif VRY > "1110000100" then--1001011000
			SY <= "10";
			s1 <= mov2;
		else
			SY <= "11";
			s1 <= mov0;
		end if;
	---Parte Servomotor con 180� de libertad
		if relogio'event and relogio = '1' then
			if VRX < "0100101100" then
				SX <= "01";
				if se�alt = "00000" then
					se�alt <= "00000";
				else
					se�alt <= se�alt - "00001";
				end if;
			elsif VRX > "1110000100" then
				SX <= "10";
				if se�alt = "10011" then
					se�alt <= "10011";
				else
					se�alt <= se�alt + "00001";
				end if;
			else 
				SX <= "11";
				se�alt <= se�alt;
			end if;
		end if;
	end process;
--Divisor de Frecuencia para selector--
	Process(clk)begin
		if clk'event and clk = '1' then
			if cont0 = 1500000 then --1000000 = 25Hz
				cont0 <= 1;
				relogio <= not relogio;
			else
				cont0 <= cont0 + 1;
			end if;
		end if;
	end process;
----Divisor de Frecuencia cont servo libre----
	Process (clk) begin
		if clk'event and clk = '1' then
			if cont = 12500 then --12500 = 2kHz
				cont <= 1;
				uhr <= not uhr;
			else
				cont <= cont + 1;
			end if;
		end if;
	end process;
---Divisor de Frecuencia cont servo con tope---
	process (clk) begin
		if clk'event and clk = '1' then
			if cont1 = 2500 then
				cont1 <= 1;
				T <= not T;
			else
				cont1 <= cont1 + 1;
			end if;
		end if;
	end process;
-----Se�ales para servo sin tope-----
	process (uhr, se�al) begin
		if uhr'event and uhr = '1' then
			se�al <= se�al + "000001";
		else 
			se�al <= se�al;---------------------------------------------------
		end if;
		case se�al is
			when "000000" =>
				mov0 <= '1';
				mov1 <= '1';
				mov2 <= '1';
			when "000001" =>
				mov0 <= '1';
				mov1 <= '1';
				mov2 <= '1';
			when "000010" =>
				mov0 <= '1';
				mov1 <= '0';
				mov2 <= '1';
			when "000011" =>
				mov0 <= '0';
				mov1 <= '0';
				mov2 <= '1';
			when "000100" =>
				mov0 <= '0';
				mov1 <= '0';
				mov2 <= '0';
			when others => 
				mov0 <= '0';
				mov1 <= '0';
				mov2 <= '0';
		end case;
	end process;
-----Se�ales para servo con tope-----
	process (se�alt,s�0,s�1,s�2,s�3,s�4,s�5,s�6,s�7,s�8,s�9,
				s�10,s�11,s�12,s�13,s�14,s�15,s�16,s�17,s�18,s�19) begin
		case se�alt is --se�alt es de 4 bits
			when "00000" => s2 <= s�0;
			when "00001" => s2 <= s�1;
			when "00010" => s2 <= s�2;
			when "00011" => s2 <= s�3;
			when "00100" => s2 <= s�4;
			when "00101" => s2 <= s�5;
			when "00110" => s2 <= s�6;
			when "00111" => s2 <= s�7;
			when "01000" => s2 <= s�8;
			when "01001" => s2 <= s�9;
			when "01010" => s2 <= s�10;
			when "01011" => s2 <= s�11;
			when "01100" => s2 <= s�12;
			when "01101" => s2 <= s�13;
			when "01110" => s2 <= s�14;
			when "01111" => s2 <= s�15;
			when "10000" => s2 <= s�16;
			when "10001" => s2 <= s�17;
			when "10010" => s2 <= s�18;
			when "10011" => s2 <= s�19;
			when others => s2 <= s�8;
		end case;
	end process;
	process (T,doscientos) begin
		if T'event and T = '1' then
			doscientos <= doscientos + "00000001";
		end if;
		case doscientos is
			when "00000000" => --1
				s�0 <= '1';
				s�1 <= '1';
				s�2 <= '1';
				s�3 <= '1';
				s�4 <= '1';
				s�5 <= '1';
				s�6 <= '1';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00000001" => --2
				s�0 <= '1';
				s�1 <= '1';
				s�2 <= '1';
				s�3 <= '1';
				s�4 <= '1';
				s�5 <= '1';
				s�6 <= '1';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00000010" => --3
				s�0 <= '1';
				s�1 <= '1';
				s�2 <= '1';
				s�3 <= '1';
				s�4 <= '1';
				s�5 <= '1';
				s�6 <= '1';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00000011" => --4
				s�0 <= '1';
				s�1 <= '1';
				s�2 <= '1';
				s�3 <= '1';
				s�4 <= '1';
				s�5 <= '1';
				s�6 <= '1';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
		---------------------------
			when "00000100" => --5
				s�0 <= '0';
				s�1 <= '1';
				s�2 <= '1';
				s�3 <= '1';
				s�4 <= '1';
				s�5 <= '1';
				s�6 <= '1';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00000101" => --6
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '1';
				s�3 <= '1';
				s�4 <= '1';
				s�5 <= '1';
				s�6 <= '1';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00000110" => --7
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '1';
				s�4 <= '1';
				s�5 <= '1';
				s�6 <= '1';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00000111" => --8
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '1';
				s�5 <= '1';
				s�6 <= '1';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00001000" => --9
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '1';
				s�6 <= '1';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00001001" => --10
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '1';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00001010" => --11
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00001011" => --12
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00001100" => --13
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00001101" => --14
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '0';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00001110" => --15
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '0';
				s�10 <= '0';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00001111" => --16
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '0';
				s�10 <= '0';
				s�11 <= '0';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00010000" => --17
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '0';
				s�10 <= '0';
				s�11 <= '0';
				s�12 <= '0';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00010001" => --18
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '0';
				s�10 <= '0';
				s�11 <= '0';
				s�12 <= '0';
				s�13 <= '0';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00010010" => --19
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '0';
				s�10 <= '0';
				s�11 <= '0';
				s�12 <= '0';
				s�13 <= '0';
				s�14 <= '0';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00010011" => --20
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '0';
				s�10 <= '0';
				s�11 <= '0';
				s�12 <= '0';
				s�13 <= '0';
				s�14 <= '0';
				s�15 <= '0';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00010100" => --21
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '0';
				s�10 <= '0';
				s�11 <= '0';
				s�12 <= '0';
				s�13 <= '0';
				s�14 <= '0';
				s�15 <= '0';
				s�16 <= '0';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when "00010101" => --22
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '0';
				s�10 <= '0';
				s�11 <= '0';
				s�12 <= '0';
				s�13 <= '0';
				s�14 <= '0';
				s�15 <= '0';
				s�16 <= '0';
				s�17 <= '0';
				s�18 <= '1';
				s�19 <= '1';
			when "00010110" => --23
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0'; 
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '0';
				s�10 <= '0';
				s�11 <= '0';
				s�12 <= '0';
				s�13 <= '0';
				s�14 <= '0';
				s�15 <= '0';
				s�16 <= '0';
				s�17 <= '0';
				s�18 <= '0';
				s�19 <= '1';
			when "11111111" => 
				s�0 <= '1';
				s�1 <= '1';
				s�2 <= '1';
				s�3 <= '1';
				s�4 <= '1';
				s�5 <= '1';
				s�6 <= '1';
				s�7 <= '1';
				s�8 <= '1';
				s�9 <= '1';
				s�10 <= '1';
				s�11 <= '1';
				s�12 <= '1';
				s�13 <= '1';
				s�14 <= '1';
				s�15 <= '1';
				s�16 <= '1';
				s�17 <= '1';
				s�18 <= '1';
				s�19 <= '1';
			when others =>
				s�0 <= '0';
				s�1 <= '0';
				s�2 <= '0';
				s�3 <= '0';
				s�4 <= '0';
				s�5 <= '0';
				s�6 <= '0';
				s�7 <= '0';
				s�8 <= '0';
				s�9 <= '0';
				s�10 <= '0';
				s�11 <= '0';
				s�12 <= '0';
				s�13 <= '0';
				s�14 <= '0';
				s�15 <= '0';
				s�16 <= '0';
				s�17 <= '0';
				s�18 <= '0';
				s�19 <= '0';
		end case;
	end process;
end Behavioral;

